interface intf();
   
    logic s;
    logic r;
    logic q;
    logic qbar;
    
        
endinterface
